** sch_path: /foss/designs/Tiny_Tapeout/TTIHP0p3_HBT_555_Timer/xschem/TB_SR_latch.sch
**.subckt TB_SR_latch
Vsrc_agnd agnd GND 0
Vsrc_avdd avdd agnd 1.8
Vsrc_S S agnd PULSE(0 1.8 0 0.5u 0.5u 3u 6u)
x1 avdd Q_bar Q agnd S R SR_latch
Vsrc_R R agnd PULSE(0 1.8 0 0.5u 0.5u 4u 8u)
x9 avdd Q Q_Buf agnd buffer
x10 avdd Q_bar Q_bar_Buf agnd buffer
**** begin user architecture code


.lib /foss/designs/IHP-Open-PDK/ihp-sg13g2/libs.tech/ngspice/models/cornerHBT.lib hbt_typ
.lib /foss/designs/IHP-Open-PDK/ihp-sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ
.lib /foss/designs/IHP-Open-PDK/ihp-sg13g2/libs.tech/ngspice/models/cornerCAP.lib cap_typ
.lib /foss/designs/IHP-Open-PDK/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt

.include /foss/designs/IHP-Open-PDK/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice

*.lib /foss/designs/IHP-Open-PDK/ihp-sg13g2/libs.tech/ngspice/models/cornerHBT.lib hbt_typ_stat
*.lib /foss/designs/IHP-Open-PDK/ihp-sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ_stat

*.lib /foss/designs/IHP-Open-PDK/ihp-sg13g2/libs.tech/ngspice/models/resistors_stat.lib
*.lib /foss/designs/IHP-Open-PDK/ihp-sg13g2/libs.tech/ngspice/models/resistors_mod.lib

* this option enables mos model bin
* selection based on W/NF instead of W
.option wnflag=1

.option savecurrents

.control
save all
op

* Print newline
echo

* Stimulus voltage
*Vstim stim 0 DC=0V
*.param Vstim = PWL(0 0 1u 1.8 2u 0 3u 1.8 4u 0)

* Sweep frequency and time
write TB_SR_latch.raw
set appendwrite

* Analyses
ac dec 100 1 1e11
tran 10n 40u
*dc vsrc_stim 0 1.8 0.1
remzerovec

* Inputs
let vin_S = v(S)
let vin_R = v(R)

* Outputs
let vout_Q = v(Q)
let vout_Q_bar = v(Q_bar)

* Plot outputs
*plot v(VB_2)
*plot v(VB_1)
*plot v(stim)

write TB_SR_latch.raw
set appendwrite

.endc


**** end user architecture code
**.ends

* expanding   symbol:  SR_latch.sym # of pins=6
** sym_path: /foss/designs/Tiny_Tapeout/TTIHP0p3_HBT_555_Timer/xschem/SR_latch.sym
** sch_path: /foss/designs/Tiny_Tapeout/TTIHP0p3_HBT_555_Timer/xschem/SR_latch.sch
.subckt SR_latch avdd Q_bar Q agnd S R
*.ipin R
*.opin Q_bar
*.ipin S
*.opin Q
*.iopin avdd
*.iopin agnd
XQ2 Q_bar net2 agnd agnd npn13G2 Nx=1
XQ1 Q net1 agnd agnd npn13G2 Nx=1
XR3 R net1 rppd w=0.5e-6 l=20e-6 m=1 b=0
XR1 net2 S rppd w=0.5e-6 l=20e-6 m=1 b=0
XR2 agnd net1 rhigh w=0.5e-6 l=20e-6 m=1 b=0
XR4 agnd net2 rhigh w=0.5e-6 l=20e-6 m=1 b=0
XR5 Q net2 rppd w=0.5e-6 l=20e-6 m=1 b=0
XR6 net1 Q_bar rppd w=0.5e-6 l=20e-6 m=1 b=0
XR7 Q avdd rppd w=0.5e-6 l=2e-6 m=1 b=0
XR8 Q_bar avdd rppd w=0.5e-6 l=2e-6 m=1 b=0
.ends


* expanding   symbol:  buffer.sym # of pins=4
** sym_path: /foss/designs/Tiny_Tapeout/TTIHP0p3_HBT_555_Timer/xschem/buffer.sym
** sch_path: /foss/designs/Tiny_Tapeout/TTIHP0p3_HBT_555_Timer/xschem/buffer.sch
.subckt buffer avdd vin vout agnd
*.iopin avdd
*.ipin vin
*.opin vout
*.iopin agnd
x1 avdd vin net1 agnd inverter
x2 avdd net1 vout agnd inverter
.ends


* expanding   symbol:  inverter.sym # of pins=4
** sym_path: /foss/designs/Tiny_Tapeout/TTIHP0p3_HBT_555_Timer/xschem/inverter.sym
** sch_path: /foss/designs/Tiny_Tapeout/TTIHP0p3_HBT_555_Timer/xschem/inverter.sch
.subckt inverter avdd vin vout agnd
*.iopin avdd
*.ipin vin
*.opin vout
*.iopin agnd
XQ1 vout base agnd agnd npn13G2 Nx=10
XR1 vout avdd rhigh w=1e-6 l=0.5e-6 m=1 b=0
XR2 vin base rhigh w=0.5e-6 l=0.5e-6 m=1 b=0
.ends

.GLOBAL GND
.end
