VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_NicklausThompson_555_1x1
  CLASS BLOCK ;
  FOREIGN tt_um_NicklausThompson_555_1x1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.000 BY 1.000 ;
END tt_um_NicklausThompson_555_1x1
END LIBRARY

