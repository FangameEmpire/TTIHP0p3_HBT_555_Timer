  X �     ,�     , LIB  >A�7KƧ�9D�/��ZT �     ,�     , tt_um_template_1x1_analog     C   ,     �d     ��  � ��  � �d     �d      C   ,     ��     �h  � �h  � ��     ��      C   ,     cd     f�  � f�  � cd     cd      C   ,     $�     (h  � (h  � $�     $�      C   ,  >�      >� U�  G U�  G      >�          C   ,  N       N  U�  V� U�  V�      N           C   , ڪ Y| ڪ ]d �� ]d �� Y| ڪ Y| +  ,clk       C   , � Y| � ]d �� ]d �� Y| � Y| +  ,ena       C   , ˪ Y| ˪ ]d �� ]d �� Y| ˪ Y| +  
,rst_n       C   , �� Y| �� ]d �� ]d �� Y| �� Y| +  ,ui_in[0]      C   , �� Y| �� ]d �� ]d �� Y| �� Y| +  ,ui_in[1]      C   , �� Y| �� ]d �� ]d �� Y| �� Y| +  ,ui_in[2]      C   , �� Y| �� ]d �� ]d �� Y| �� Y| +  ,ui_in[3]      C   , �� Y| �� ]d �� ]d �� Y| �� Y| +  ,ui_in[4]      C   , q� Y| q� ]d r� ]d r� Y| q� Y| +  ,ui_in[5]      C   , b� Y| b� ]d c� ]d c� Y| b� Y| +  ,ui_in[6]      C   , S� Y| S� ]d T� ]d T� Y| S� Y| +  ,ui_in[7]      C   , D� Y| D� ]d E� ]d E� Y| D� Y| +  ,uio_in[0]       C   , 5� Y| 5� ]d 6� ]d 6� Y| 5� Y| +  ,uio_in[1]       C   , &� Y| &� ]d '� ]d '� Y| &� Y| +  ,uio_in[2]       C   , � Y| � ]d � ]d � Y| � Y| +  ,uio_in[3]       C   , � Y| � ]d 	� ]d 	� Y| � Y| +  ,uio_in[4]       C   , �� Y| �� ]d �� ]d �� Y| �� Y| +  ,uio_in[5]       C   , � Y| � ]d �� ]d �� Y| � Y| +  ,uio_in[6]       C   , ۪ Y| ۪ ]d �� ]d �� Y| ۪ Y| +  ,uio_in[7]       C   ,  ܪ Y|  ܪ ]d  �� ]d  �� Y|  ܪ Y| +  ,uio_oe[0]       C   ,  ͪ Y|  ͪ ]d  �� ]d  �� Y|  ͪ Y| +  ,uio_oe[1]       C   ,  �� Y|  �� ]d  �� ]d  �� Y|  �� Y| +  ,uio_oe[2]       C   ,  �� Y|  �� ]d  �� ]d  �� Y|  �� Y| +  ,uio_oe[3]       C   ,  �� Y|  �� ]d  �� ]d  �� Y|  �� Y| +  ,uio_oe[4]       C   ,  �� Y|  �� ]d  �� ]d  �� Y|  �� Y| +  ,uio_oe[5]       C   ,  �� Y|  �� ]d  �� ]d  �� Y|  �� Y| +  ,uio_oe[6]       C   ,  s� Y|  s� ]d  t� ]d  t� Y|  s� Y| +  ,uio_oe[7]       C   , T� Y| T� ]d U� ]d U� Y| T� Y| +  ,uio_out[0]      C   , E� Y| E� ]d F� ]d F� Y| E� Y| +  ,uio_out[1]      C   , 6� Y| 6� ]d 7� ]d 7� Y| 6� Y| +  ,uio_out[2]      C   , '� Y| '� ]d (� ]d (� Y| '� Y| +  ,uio_out[3]      C   , � Y| � ]d � ]d � Y| � Y| +  ,uio_out[4]      C   , 	� Y| 	� ]d 
� ]d 
� Y| 	� Y| +  ,uio_out[5]      C   ,  �� Y|  �� ]d  �� ]d  �� Y|  �� Y| +  ,uio_out[6]      C   ,  � Y|  � ]d  �� ]d  �� Y|  � Y| +  ,uio_out[7]      C   , ̪ Y| ̪ ]d �� ]d �� Y| ̪ Y| +  ,uo_out[0]       C   , �� Y| �� ]d �� ]d �� Y| �� Y| +  ,uo_out[1]       C   , �� Y| �� ]d �� ]d �� Y| �� Y| +  ,uo_out[2]       C   , �� Y| �� ]d �� ]d �� Y| �� Y| +  ,uo_out[3]       C   , �� Y| �� ]d �� ]d �� Y| �� Y| +  ,uo_out[4]       C   , �� Y| �� ]d �� ]d �� Y| �� Y| +  ,uo_out[5]       C   , r� Y| r� ]d s� ]d s� Y| r� Y| +  ,uo_out[6]       C   , c� Y| c� ]d d� ]d d� Y| c� Y| +  ,uo_out[7]       �   ,             ]d ` ]d `                  C    , ڪ Y| ڪ ]d �� ]d �� Y| ڪ Y|      C    , � Y| � ]d �� ]d �� Y| � Y|      C    , ˪ Y| ˪ ]d �� ]d �� Y| ˪ Y|      C    , �� Y| �� ]d �� ]d �� Y| �� Y|      C    , �� Y| �� ]d �� ]d �� Y| �� Y|      C    , �� Y| �� ]d �� ]d �� Y| �� Y|      C    , �� Y| �� ]d �� ]d �� Y| �� Y|      C    , �� Y| �� ]d �� ]d �� Y| �� Y|      C    , q� Y| q� ]d r� ]d r� Y| q� Y|      C    , b� Y| b� ]d c� ]d c� Y| b� Y|      C    , S� Y| S� ]d T� ]d T� Y| S� Y|      C    , D� Y| D� ]d E� ]d E� Y| D� Y|      C    , 5� Y| 5� ]d 6� ]d 6� Y| 5� Y|      C    , &� Y| &� ]d '� ]d '� Y| &� Y|      C    , � Y| � ]d � ]d � Y| � Y|      C    , � Y| � ]d 	� ]d 	� Y| � Y|      C    , �� Y| �� ]d �� ]d �� Y| �� Y|      C    , � Y| � ]d �� ]d �� Y| � Y|      C    , ۪ Y| ۪ ]d �� ]d �� Y| ۪ Y|      C    ,  ܪ Y|  ܪ ]d  �� ]d  �� Y|  ܪ Y|      C    ,  ͪ Y|  ͪ ]d  �� ]d  �� Y|  ͪ Y|      C    ,  �� Y|  �� ]d  �� ]d  �� Y|  �� Y|      C    ,  �� Y|  �� ]d  �� ]d  �� Y|  �� Y|      C    ,  �� Y|  �� ]d  �� ]d  �� Y|  �� Y|      C    ,  �� Y|  �� ]d  �� ]d  �� Y|  �� Y|      C    ,  �� Y|  �� ]d  �� ]d  �� Y|  �� Y|      C    ,  s� Y|  s� ]d  t� ]d  t� Y|  s� Y|      C    , T� Y| T� ]d U� ]d U� Y| T� Y|      C    , E� Y| E� ]d F� ]d F� Y| E� Y|      C    , 6� Y| 6� ]d 7� ]d 7� Y| 6� Y|      C    , '� Y| '� ]d (� ]d (� Y| '� Y|      C    , � Y| � ]d � ]d � Y| � Y|      C    , 	� Y| 	� ]d 
� ]d 
� Y| 	� Y|      C    ,  �� Y|  �� ]d  �� ]d  �� Y|  �� Y|      C    ,  � Y|  � ]d  �� ]d  �� Y|  � Y|      C    , ̪ Y| ̪ ]d �� ]d �� Y| ̪ Y|      C    , �� Y| �� ]d �� ]d �� Y| �� Y|      C    , �� Y| �� ]d �� ]d �� Y| �� Y|      C    , �� Y| �� ]d �� ]d �� Y| �� Y|      C    , �� Y| �� ]d �� ]d �� Y| �� Y|      C    , �� Y| �� ]d �� ]d �� Y| �� Y|      C    , r� Y| r� ]d s� ]d s� Y| r� Y|      C    , c� Y| c� ]d d� ]d d� Y| c� Y|      C    ,     �d     ��  � ��  � �d     �d      C    ,     ��     �h  � �h  � ��     ��      C    ,     cd     f�  � f�  � cd     cd      C    ,     $�     (h  � (h  � $�     $�      C    ,  >�      >� U�  G U�  G      >�          C    ,  N       N  U�  V� U�  V�      N           C       �@ [p clk       C       �@ [p ena       C       �@ [p 
rst_n       C       �@ [p ui_in[0]      C       �@ [p ui_in[1]      C       �@ [p ui_in[2]      C       �@ [p ui_in[3]      C       �@ [p ui_in[4]      C       r@ [p ui_in[5]      C       c@ [p ui_in[6]      C       T@ [p ui_in[7]      C       E@ [p uio_in[0]       C       6@ [p uio_in[1]       C       '@ [p uio_in[2]       C       @ [p uio_in[3]       C       	@ [p uio_in[4]       C       �@ [p uio_in[5]       C       �@ [p uio_in[6]       C       �@ [p uio_in[7]       C        �@ [p uio_oe[0]       C        �@ [p uio_oe[1]       C        �@ [p uio_oe[2]       C        �@ [p uio_oe[3]       C        �@ [p uio_oe[4]       C        �@ [p uio_oe[5]       C        �@ [p uio_oe[6]       C        t@ [p uio_oe[7]       C       U@ [p uio_out[0]      C       F@ [p uio_out[1]      C       7@ [p uio_out[2]      C       (@ [p uio_out[3]      C       @ [p uio_out[4]      C       
@ [p uio_out[5]      C        �@ [p uio_out[6]      C        �@ [p uio_out[7]      C       �@ [p uo_out[0]       C       �@ [p uo_out[1]       C       �@ [p uo_out[2]       C       �@ [p uo_out[3]       C       �@ [p uo_out[4]       C       �@ [p uo_out[5]       C       s@ [p uo_out[6]       C       d@ [p uo_out[7]       C       � �& 
ua[0]       C       � �� 
ua[1]       C       � e& 
ua[2]       C       � &� 
ua[3]       C       B� *� VGND      C       Rl *� VPWR      