** sch_path: /foss/designs/Tiny_Tapeout/TTIHP0p3_HBT_555_Timer/xschem/TB_555.sch
**.subckt TB_555
x1 avdd VB_1 555_Vout VB_2 VB_1 agnd 555
Vsrc_agnd agnd GND 0
Vsrc_avdd avdd agnd 1.8
C1 VB_1 agnd 10n m=1
R1 avdd VB_2 1k m=1
R2 VB_2 VB_1 1k m=1
**** begin user architecture code


.lib /foss/designs/IHP-Open-PDK/ihp-sg13g2/libs.tech/ngspice/models/cornerHBT.lib hbt_typ
.lib /foss/designs/IHP-Open-PDK/ihp-sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ
.lib /foss/designs/IHP-Open-PDK/ihp-sg13g2/libs.tech/ngspice/models/cornerCAP.lib cap_typ
.lib /foss/designs/IHP-Open-PDK/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt

.include /foss/designs/IHP-Open-PDK/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice

*.lib /foss/designs/IHP-Open-PDK/ihp-sg13g2/libs.tech/ngspice/models/cornerHBT.lib hbt_typ_stat
*.lib /foss/designs/IHP-Open-PDK/ihp-sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ_stat

*.lib /foss/designs/IHP-Open-PDK/ihp-sg13g2/libs.tech/ngspice/models/resistors_stat.lib
*.lib /foss/designs/IHP-Open-PDK/ihp-sg13g2/libs.tech/ngspice/models/resistors_mod.lib

* this option enables mos model bin
* selection based on W/NF instead of W
.option wnflag=1

.option savecurrents

.control
save all
op

* Print newline
echo

* Analyses
tran 0.1u 400u
remzerovec

* Inputs


* Outputs


* Plot outputs


write TB_555.raw
set appendwrite

.endc


**** end user architecture code
**.ends

* expanding   symbol:  555.sym # of pins=6
** sym_path: /foss/designs/Tiny_Tapeout/TTIHP0p3_HBT_555_Timer/xschem/555.sym
** sch_path: /foss/designs/Tiny_Tapeout/TTIHP0p3_HBT_555_Timer/xschem/555.sch
.subckt 555 avdd THRESHOLD OUT DISCHARGE TRIGGER agnd
*.opin OUT
*.iopin avdd
*.iopin agnd
*.iopin TRIGGER
*.iopin THRESHOLD
*.iopin DISCHARGE
XR3 VB_2 avdd rhigh w=0.5e-6 l=1.59e-6 m=1 b=0
XR1 agnd VB_1 rhigh w=0.5e-6 l=1.59e-6 m=1 b=0
XR2 VB_1 VB_2 rhigh w=0.5e-6 l=1.59e-6 m=1 b=0
XC1 VB_1 agnd cap_cmim w=7.0e-6 l=7.0e-6 m=1
XC2 VB_2 agnd cap_cmim w=7.0e-6 l=7.0e-6 m=1
XC3 avdd agnd cap_cmim w=7.0e-6 l=7.0e-6 m=1
XR4 out_bar net7 rhigh w=0.5e-6 l=1.59e-6 m=1 b=0
x1 avdd net2 net8 VB_2 THRESHOLD agnd comparator
x2 avdd net1 net9 TRIGGER VB_1 agnd comparator
x9 avdd net2 net4 agnd buffer
x10 avdd net1 net3 agnd buffer
x3 avdd net6 net5 agnd net3 net4 SR_latch
x4 avdd net5 OUT agnd buffer
x5 avdd net6 out_bar agnd buffer
* noconn #net8
* noconn #net9
XQ1 DISCHARGE net7 agnd agnd npn13G2 Nx=1
.ends


* expanding   symbol:  comparator.sym # of pins=6
** sym_path: /foss/designs/Tiny_Tapeout/TTIHP0p3_HBT_555_Timer/xschem/comparator.sym
** sch_path: /foss/designs/Tiny_Tapeout/TTIHP0p3_HBT_555_Timer/xschem/comparator.sch
.subckt comparator avdd voutp voutn vinn vinp agnd
*.iopin avdd
*.ipin vinp
*.opin voutp
*.iopin agnd
*.ipin vinn
*.opin voutn
XQ1 voutp vinn ee agnd npn13G2 Nx=1
XR1 voutp avdd rppd w=0.5e-6 l=30e-6 m=1 b=0
XR2 agnd ee rppd w=0.5e-6 l=0.5e-6 m=1 b=0
XR3 voutn avdd rppd w=0.5e-6 l=30e-6 m=1 b=0
XQ2 voutn vinp ee agnd npn13G2 Nx=1
.ends


* expanding   symbol:  buffer.sym # of pins=4
** sym_path: /foss/designs/Tiny_Tapeout/TTIHP0p3_HBT_555_Timer/xschem/buffer.sym
** sch_path: /foss/designs/Tiny_Tapeout/TTIHP0p3_HBT_555_Timer/xschem/buffer.sch
.subckt buffer avdd vin vout agnd
*.iopin avdd
*.ipin vin
*.opin vout
*.iopin agnd
x1 avdd vin net1 agnd inverter
x2 avdd net1 vout agnd inverter
.ends


* expanding   symbol:  SR_latch.sym # of pins=6
** sym_path: /foss/designs/Tiny_Tapeout/TTIHP0p3_HBT_555_Timer/xschem/SR_latch.sym
** sch_path: /foss/designs/Tiny_Tapeout/TTIHP0p3_HBT_555_Timer/xschem/SR_latch.sch
.subckt SR_latch avdd Q_bar Q agnd S R
*.ipin R
*.opin Q_bar
*.ipin S
*.opin Q
*.iopin avdd
*.iopin agnd
XQ2 Q_bar net2 agnd agnd npn13G2 Nx=1
XQ1 Q net1 agnd agnd npn13G2 Nx=1
XR3 R net1 rppd w=0.5e-6 l=20e-6 m=1 b=0
XR1 net2 S rppd w=0.5e-6 l=20e-6 m=1 b=0
XR2 agnd net1 rhigh w=0.5e-6 l=20e-6 m=1 b=0
XR4 agnd net2 rhigh w=0.5e-6 l=20e-6 m=1 b=0
XR5 Q net2 rppd w=0.5e-6 l=20e-6 m=1 b=0
XR6 net1 Q_bar rppd w=0.5e-6 l=20e-6 m=1 b=0
XR7 Q avdd rppd w=0.5e-6 l=2e-6 m=1 b=0
XR8 Q_bar avdd rppd w=0.5e-6 l=2e-6 m=1 b=0
.ends


* expanding   symbol:  inverter.sym # of pins=4
** sym_path: /foss/designs/Tiny_Tapeout/TTIHP0p3_HBT_555_Timer/xschem/inverter.sym
** sch_path: /foss/designs/Tiny_Tapeout/TTIHP0p3_HBT_555_Timer/xschem/inverter.sch
.subckt inverter avdd vin vout agnd
*.iopin avdd
*.ipin vin
*.opin vout
*.iopin agnd
XQ1 vout base agnd agnd npn13G2 Nx=10
XR1 vout avdd rhigh w=1e-6 l=0.5e-6 m=1 b=0
XR2 vin base rhigh w=0.5e-6 l=0.5e-6 m=1 b=0
.ends

.GLOBAL GND
.end
